`timescale 1ns / 1ps
`include "interfaces.vh"
// URAM-to-Event buffer.
// This interfaces with pueo_uram_v3+ only!
//
// We don't need a memclk_sync here -
// pueo_uram_v3+ syncs up the readout requests
// to a phase, so begin_i always occurs in phase 1.
// It's the critical timing element.
//
// The goal here is to produce an output stream
// to feed into DOUT: we only need to output 1
// every 2 clocks, but the COBS encoding will
// end up buffering it anyway.
// With COBS the overhead is (n/254) rounded up, max:
// our data is 12,288 bytes meaning we'll pick up
// at most 49 bytes overhead. With 8 buffers that's
// 392 bytes at most. We also have the
// header as well, which is probably just going to be
//
// <event number> 4 bytes
// <event clock> 4 bytes
// so that's an additional 64 total bytes.
// Smallest FIFO we have is a single FIFO18
// which is 8x2048 so this isn't a problem.
//
// NOTE: rst_i is in memclk domain
//       ifclk_rst_i is in ifclk domain
//       Resets here need to be applied
//       -> assert ifclk reset
//       -> assert memclk reset
//       -> release memclk reset
//       -> release ifclk reset
//       and the resets obviously need to be held for a minimum # of clocks (16 is good enough for all of ours)
// We need an overall reset controller which sequences stuff. Our overall goal is to
// keep the reset inputs at each module as simple as possible and allow them to be pipelined.

// We also now generate an event header as well,
// containing a 2-byte event number and the 2-byte
// trigger time.
// We have a very small buffer here (16 entries, using
// distram) to hold the trigger time. Because the read
// into the event buffer takes macroscopic time (342 ns)
// there's no worry here, it will always be ready first.
//
// The annoying thing here is that it means we now need
// to register the final output to mux it, and we also have
// to wait for the data to finish outputting before we totally complete.
// WHATEVER.
//
// NOTE NOTE NOTE NOTE NOTE NOTE NOTE
// This module produces valid new data when syncclk_phase is HIGH
// tvalid is asserted then.
module uram_event_buffer #(parameter NCHAN = 8,
                           parameter NBIT_IN = 72,
                           parameter BEGIN_PHASE = 1,
                           parameter DOUT_LATENCY = 6)(
        input memclk_i,
        input memclk_rst_i,
        input begin_i,
        input [NBIT_IN*NCHAN-1:0] dat_i,
        input [NCHAN-1:0] dat_valid_i,
        input ifclk_rst_i,
        output write_error_o,
        // the input here just becomes valid every
        // other clock until the last
        input ifclk_i,
        // trigger time input
        input [14:0] trig_time_i,
        input [15:0] event_no_i,
        input        trig_valid_i,
        // fw update stuff
        input [7:0]  fw_dat_i,
        input        fw_wr_i,
        // comes from idctrl
        input        fw_load_i,
        // output data. 
        output [7:0] dout_data_o,
        output       dout_data_valid_o,
        output       dout_data_last_o,
        input        dout_data_phase_i
    );
    
    // whatever!! I'll figure out write error later
    // or maybe never at all
    assign write_error_o = 1'b0;
    
    // NOTE: BEGIN_DELAY needs to be structured so that the address arrives
    // *** 1 AFTER *** THE DATA
    // THE DATA IS GOING TO BE DELAYED BY THE MUX/REREGISTER    
    localparam BEGIN_DELAY = 6;
    localparam [3:0] BEGIN_DELAY_VAL = (BEGIN_DELAY == 0) ? 0 : BEGIN_DELAY-1;
    wire begin_delayed;
    wire this_begin = (BEGIN_DELAY == 0) ? begin_i : begin_delayed;
    SRL16E u_begin_delay(.D(begin_i),
                         .CE(1'b1),
                         .CLK(memclk_i),
                         .A0(BEGIN_DELAY_VAL[0]),
                         .A1(BEGIN_DELAY_VAL[1]),
                         .A2(BEGIN_DELAY_VAL[2]),
                         .A3(BEGIN_DELAY_VAL[3]),
                         .Q(begin_delayed));
    
    // The details here are documented in the event buffer section
    // of the firmware documentation.
    // This is trickier than it first seems.
    
    // Nominally we start off by cascading the entire thing:
    // 24 total block RAMs (8 ch x 3 per channel).
    // Writing occurs at memclk speed (500 MHz), reading at ifclk speed (125 MHz)
    // So writing needs to be easy.
    
    // We write 3 addresses (24 samples) per 4 clock cycles.
    // We will ALWAYS get begin_i in phase 1.
    // Let's just consider channel 0 for the moment.
    // Suppose we register begin_i: this will then go high in phase 2.
    // We then use this signal to reset the address generation, so it's reset in phase 3.
    // The timing of a 4-address increment will always be
    // 5/6/5 6/5/6
    // This pattern is generated by the uram_event_timer.
    // We generate a global next upper address which gets captured by ch0 and
    // forwarded.
    wire [7:0] next_bram_uaddr[NCHAN-1:0];
    // the top 3 bits are the buffer. They're Gray encoded so they can
    // hop across domains. Thankfully a 3-bit Gray counter fits in logic.

    // This is the *in progress* buffer pointer.
    // This gets incremented when the first channel finishes.
    reg [2:0] write_buffer = {3{1'b0}};
    // This is the *completed* buffer pointer. This gets incremented
    // when the last channel finishes.
    reg [2:0] complete_buffer_pointer = {3{1'b0}};
    // The reason we have 2 buffer pointers is because our control logic
    // is pipelined. We could probably just start reading out early,
    // but I'd rather be safe than sorry.
    
    // This is the upper address pointer.
    // We only pass the top 5 bits to the individual channels.
    reg [4:0] write_addr = {5{1'b0}};    
    reg [1:0] glob_memclk_phase = {2{1'b0}};
    localparam [1:0] GLOB_MEMCLK_PHASE_RESET_VAL = 3;
    wire glob_start;
    reg running = 0;
    wire increment_uaddr;
    uram_event_timer u_timer(.memclk_i(memclk_i),
                             .memclk_phase_i(!glob_memclk_phase[0]),
                             .running_i(running),
                             .start_o(glob_start),
                             .capture_o(increment_uaddr));
    // ok we still need to figure out when to *terminate* running
    localparam TERMINATE_VAL = {5{1'b1}};
    // and then once we hit that point, we need
    // to delay the terminate slightly to line everything
    // up. The URAM reads out 1026 samples: looking at the
    // physical transition flow you can see that it'll
    // be phase 3 that we stop at, because the 'stored'
    // A0/A1/A2 data (2 samples) will be discarded.
    // If you work out the logic you'd *expect* this to be 2
    // but the extra clock comes because we don't increment
    // in phase 1.
    //
    // Working it out, after this_begin goes high,
    // the next this_begin cannot occur for another 350 ns,
    // or 175 clocks: in other words, we add *one* 4-clock
    // period for every event we're actively reading out.
    //
    // We can probably just integrate this timing into the trigger
    // readout at the TURF since everything's synchronous.
    localparam TERMINATE_DELAY = 3;    
    localparam [3:0] SRL_TERMINATE_DELAY = TERMINATE_DELAY-1;
    reg terminate_seen = 0;
    wire do_terminate;
    // we use terminate_seen to act as a portion of our
    // reset - but that means it needs to be a flag
    reg memclk_reset = 0;
    reg memclk_reset_rereg = 0;
    reg memclk_reset_flag = 0;
    
    SRL16E u_terminate_delay(.D(terminate_seen),
                             .CE(1'b1),
                             .CLK(memclk_i),
                             .A0(SRL_TERMINATE_DELAY[0]),
                             .A1(SRL_TERMINATE_DELAY[1]),
                             .A2(SRL_TERMINATE_DELAY[2]),
                             .A3(SRL_TERMINATE_DELAY[3]),
                             .Q(do_terminate));
    // and then we also need to have a complete delay
    // to signal the other side that we have an event
    // ready to read out.
    localparam COMPLETE_DELAY = 31;
    localparam [4:0] SRL_COMPLETE_DELAY = COMPLETE_DELAY-1;
    wire do_complete;
    SRLC32E u_complete_delay(.D(do_terminate),
                             .CE(1'b1),
                             .CLK(memclk_i),
                             .A(SRL_COMPLETE_DELAY),
                             .Q(do_complete));
                                 
    always @(posedge memclk_i) begin
        memclk_reset <= memclk_rst_i;
        memclk_reset_rereg <= memclk_reset;
        memclk_reset_flag <= memclk_reset && !memclk_reset_rereg;
    
        if (begin_delayed) running <= 1;
        else if (do_terminate) running <= 0;
        
        // Gray coded write buffer.
        if (memclk_reset) write_buffer <= {3{1'b0}};
        else if (do_terminate) begin
            case (write_buffer)
                3'b000: write_buffer <= 3'b001;
                3'b001: write_buffer <= 3'b011;
                3'b011: write_buffer <= 3'b010;
                3'b010: write_buffer <= 3'b110;
                3'b110: write_buffer <= 3'b111;
                3'b111: write_buffer <= 3'b101;
                3'b101: write_buffer <= 3'b100;
                3'b100: write_buffer <= 3'b000;
            endcase
        end        
        // Gray coded complete buffer pointer.
        if (memclk_reset) complete_buffer_pointer <= 3'b000;
        else if (do_complete) begin
            case (complete_buffer_pointer)
                3'b000: complete_buffer_pointer <= 3'b001;
                3'b001: complete_buffer_pointer <= 3'b011;
                3'b011: complete_buffer_pointer <= 3'b010;
                3'b010: complete_buffer_pointer <= 3'b110;
                3'b110: complete_buffer_pointer <= 3'b111;
                3'b111: complete_buffer_pointer <= 3'b101;
                3'b101: complete_buffer_pointer <= 3'b100;
                3'b100: complete_buffer_pointer <= 3'b000;
            endcase                
        end
        
        // terminate_seen going high will kill running after a small number of clocks
        // running going low will end the readout, and everything
        // resets straight away at the next start.
        terminate_seen <= ((write_addr == TERMINATE_VAL) && increment_uaddr) || memclk_reset_flag;

        if (memclk_reset) write_addr <= {5{1'b0}};
        else if (increment_uaddr) write_addr <= write_addr + 1;
        
        if (glob_start) glob_memclk_phase <= GLOB_MEMCLK_PHASE_RESET_VAL;
        else glob_memclk_phase <= glob_memclk_phase + 1;        
    end                                  

    // READOUT PROCESS
    // Even though the readout process is basically stateful
    // it's easier to treat it as something closer to a
    // FIFO, except we don't even worry about the problem of
    // overflow because the TURF protects us from it.
    // So all we need to do is recapture the complete_buffer_pointer
    // and compare it to the read_buffer_pointer, and if they're
    // not equal, we start the readout process.
    //
    // The TURF protects from overflow by keeping its *own*
    // pointers regarding received and sent triggers.
    // This makes this a little less efficient than it could be
    // but whatever.

    // current read buffer
    reg [2:0] read_buffer = {3{1'b0}};
    // write buffer in read domain
    reg [2:0] completed_ifclk_sync = {3{1'b0}};
    // actual version to use
    reg [2:0] completed_buffer = {3{1'b0}};
    
    // once we have a buffer to read, the sequence basically looks like
    // en   addr    casdomux_i  casdomuxen_i    dout
    // 000  003     24'hFFFFFE  0               X
    // 001  000     24'hFFFFFE  1               X
    // 001  001     24'hFFFFFC  0               X
    // 001  002     ..          0               ARAM[0]
    // 001  003     ..          0               ARAM[1]
    // 010  000     24'hFFFFFC  1               ARAM[2]
    // 010  001     24'hFFFFFC  0               ARAM[3]
    // etc.
    // Note that casdomux_i[1:0] actually go to bram_casdomux_i
    // but casdomux[2] actually goes to casoregimux (same with the _en).
    // because the C BRAM feeds into its pipeline register before
    // going to the next channel.
    //
    // because of the 2 clock phase the sequence actually only
    // toggles stuff every other phase.
    // the other thing to consider is the *order* to read out
    // in. Reading out bottom to top means a longer initial
    // latency but it just means a channel switch is a delay
    // to let the other data clear through.
    reg [NCHAN-1:0] bram_regce = {NCHAN{1'b0}};
    // the bram CAS and enable stuff need to cycle when
    // they're active.
    reg [2:0] active_bram = 3'b001;
    wire [2:0] active_bram_casdomux =
        { !active_bram[2],
          !active_bram[1],
          !active_bram[0] };
    reg [NCHAN-1:0] active_chan = 8'b00000001;    
    wire [3*NCHAN-1:0] full_casdomux = {
        !active_chan[7] ? 3'b111 : active_bram_casdomux,
        !active_chan[6] ? 3'b111 : active_bram_casdomux,
        !active_chan[5] ? 3'b111 : active_bram_casdomux,
        !active_chan[4] ? 3'b111 : active_bram_casdomux,
        !active_chan[3] ? 3'b111 : active_bram_casdomux,
        !active_chan[2] ? 3'b111 : active_bram_casdomux,
        !active_chan[1] ? 3'b111 : active_bram_casdomux,
        active_bram_casdomux };
              
    reg bram_casdomuxen = 1'b0;
    // 2 address bits here. 3 for the buffer, means...
    reg [1:0] bram_lraddr = {2{1'b0}};
    // need 7 bits here
    reg [6:0] bram_uraddr = {7{1'b0}};
    wire [9:0] bram_addr = { read_buffer, bram_lraddr, bram_uraddr };
    
    // reading we can do in a state machine
    localparam FSM_BITS = 3;
    localparam [FSM_BITS-1:0] IDLE = 0;
    localparam [FSM_BITS-1:0] RESET_ALL = 1;
    localparam [FSM_BITS-1:0] CH_ADVANCE = 2;
    localparam [FSM_BITS-1:0] READING = 3;
    localparam [FSM_BITS-1:0] COMPLETE = 4;
    localparam [FSM_BITS-1:0] FW_LOAD = 5;
    reg [FSM_BITS-1:0] state = IDLE;
    reg channel_complete = 0;
    reg data_available = 0;
    reg read_terminate = 0;
    (* CUSTOM_CC_DST = "IFCLK" *)
    reg [1:0] loading_fw = {2{1'b0}};

    wire data_start = (state == RESET_ALL && dout_data_phase_i && !loading_fw[1]);
    wire data_start_delayed;
    // number of header bytes
    localparam NUM_HEADERS = 4;
    // delay from data_start to transition on event start
    // 17 clocks from data_start is when the first valid data pops
    // on last_data. The odd number is because the first bit in
    // the SRL goes high in !ifclk_phase_i: so to get a single
    // ifclk_phase delay the SRL input would need to be 1.
    localparam DATA_START_DELAY = 17 - NUM_HEADERS*2;
    localparam [4:0] SRL_VALID_DELAY_VAL = DATA_START_DELAY;
    SRLC32E u_valid_delay(.D(data_start),
                          .A(SRL_VALID_DELAY_VAL),
                          .Q(data_start_delayed),
                          .CLK(ifclk_i),
                          .CE(1'b1));
    // go high when channel_complete and active_chan[7] and !ifclk_phase_i
    reg data_tlast = 0;                          
//    // go high at data_start_delayed and go low at last                              
//    reg data_tvalid = 0;
    
    // Note: ifclk_rst_i is just treated straight since it's
    // in a slower clock domain. This means that functionally
    // its reset needs to generate the memclk reset and stay
    // in reset through.
    // Because the uram needs to handle the reset as well
    // (to terminate its reading) we generate that reset
    // sequence outside of here.
    //
    // HOW THE SLEAZEBALL WORKS
    // OUR FIRST ATTEMPT JUST USES ONE SINGLE BLOCK RAM AS A BUFFER
    // 

    always @(posedge ifclk_i) begin
        loading_fw <= { loading_fw[0], fw_load_i };
        
        if (ifclk_rst_i)
            data_tlast <= 1'b0;
        else if (!dout_data_phase_i)
            data_tlast <= channel_complete && active_chan[7];

//        if ((data_tlast && ifclk_phase_i) || ifclk_rst_i) data_tvalid <= 0;
//        else if (data_start_delayed) data_tvalid <= 1;
        
        completed_ifclk_sync <= complete_buffer_pointer;
        completed_buffer <= completed_ifclk_sync;
        data_available <= (completed_buffer != read_buffer);
        channel_complete <= ({bram_uraddr, bram_lraddr} == 9'h1FF) && active_bram[2];        
        if (state == COMPLETE || ifclk_rst_i)
            read_terminate <= 0;
        else if (channel_complete && active_chan[7])
            read_terminate <= 1;

        // this ONLY WORKS because we've got a 2-clock period
        // clk  ifclk_phase state       read_terminate read_buffer data_available
        // 0    1           CH_ADVANCE  1              0           1
        // 1    0           COMPLETE    1              0           1
        // 2    1           COMPLETE    0              1           1
        // 3    0           IDLE        0              1           0        
        if (ifclk_rst_i) read_buffer <= 3'b000;
        else if (state == COMPLETE && !dout_data_phase_i) begin
            case (read_buffer)
                3'b000: read_buffer <= 3'b001;
                3'b001: read_buffer <= 3'b011;
                3'b011: read_buffer <= 3'b010;
                3'b010: read_buffer <= 3'b110;
                3'b110: read_buffer <= 3'b111;
                3'b111: read_buffer <= 3'b101;
                3'b101: read_buffer <= 3'b100;
                3'b100: read_buffer <= 3'b000;
            endcase
        end                       

        if (ifclk_rst_i) state <= IDLE;                        
        else if (dout_data_phase_i || loading_fw[1]) begin
            case (state)
                IDLE: if (data_available || loading_fw[1]) state <= RESET_ALL;
                RESET_ALL: if (loading_fw[1]) state <= FW_LOAD;
                           else state <= CH_ADVANCE;
                CH_ADVANCE: if (read_terminate) state <= COMPLETE;
                            else state <= READING;
                READING: if (channel_complete) state <= CH_ADVANCE;               
                COMPLETE: state <= IDLE;
                FW_LOAD: if (!loading_fw[1]) state <= IDLE;
            endcase
        end
        // the weird "start with 7 and loop around" bit
        // allows us to put CH_ADVANCE in the reset process
        if (state == RESET_ALL) begin
            // hackhack. we might not need this, maybe we just
            // shove it into the top BRAM
            if (!loading_fw[1]) active_chan <= 8'b10000000;
            else active_chan <= 8'b00000001;
        end else if (state == CH_ADVANCE && dout_data_phase_i)
            active_chan <= {active_chan[6:0],active_chan[7]};

        // SIMPLE SLEAZEBALLS: EVERY TIME WE SEE A WRITE, INCREMENT
        // IT'S YOUR DAMN JOB TO FIX IT BY RESETTING
        // RIGHT NOW WITH THIS METHOD WE CAN ONLY STORE 1 BRAM WORTH
        // OF DATA 
        if (state == RESET_ALL) begin
            bram_lraddr <= 2'b00;
        end else if ((state == READING && !dout_data_phase_i) || fw_wr_i ) begin
            bram_lraddr <= bram_lraddr + 1;
        end
        if (state == RESET_ALL) begin
            active_bram <= 3'b001;
        end else if ((state == READING && !dout_data_phase_i) && bram_lraddr == 2'b11) begin
            active_bram <= {active_bram[1:0],active_bram[2]};
        end            
        if (state == RESET_ALL) begin
            bram_uraddr <= {5{1'b0}};
        end else if (((state == READING && !dout_data_phase_i && active_bram[2]) || fw_wr_i) && bram_lraddr == 2'b11) begin
            bram_uraddr <= bram_uraddr + 1;
        end            
        if (state == CH_ADVANCE) bram_casdomuxen <= 1;
        else if (state == READING && !dout_data_phase_i && bram_lraddr == 2'b11) bram_casdomuxen <= 1;
        else bram_casdomuxen <= 0;
    end

    // cascades
    wire [35:0] cas_doutb[NCHAN-1:0];
    wire [35:0] cas_dinb[NCHAN-1:0];

    assign cas_dinb[0] = {36{1'b0}};
        
    wire [7:0] last_data;
    reg [7:0]  last_data_store = {8{1'b0}};
    
    assign next_bram_uaddr[0] = { write_buffer, write_addr };
    generate
        genvar i;
        for (i=0;i<NCHAN;i=i+1) begin : CH
            wire [71:0] this_channel_data = dat_i[NBIT_IN*i +: NBIT_IN];
            wire [7:0] this_bram_uaddr = next_bram_uaddr[i];
            wire [7:0] this_next_bram_uaddr;
            
            wire [2:0] this_bram_casdomux = full_casdomux[3*i +: 3];
            wire [2:0] this_bram_casdomuxen = {3{bram_casdomuxen}};
            wire [2:0] this_bram_en = active_chan[i] ? active_bram : 3'b000;
            wire this_bram_regce = !dout_data_phase_i;
            wire [11:0] this_bram_raddr = { read_buffer, bram_uraddr, bram_lraddr };
            wire [7:0] this_bram_dat_o;
            wire [7:0] this_bram_upd_dat = {8{1'b0}};
            wire this_bram_upd_wr = 1'b0;
            wire [2:0] this_bram_upd_casdimux = {3{1'b0}};
                        
            if (i != NCHAN-1) begin : NL
                assign next_bram_uaddr[i+1] = this_next_bram_uaddr;
            end else begin
                assign last_data = this_bram_dat_o;
            end
            if (i != 0) begin : CNF
                assign cas_dinb[i] = cas_doutb[i-1];
            end
            localparam CHANNEL_ORDER = ( (i==0) ? "FIRST" : ( (i==NCHAN-1) ? "LAST" : "MIDDLE"));
            uram_event_chbuffer #(.RUN_DELAY(4*i),
                                  .CHANNEL_ORDER(CHANNEL_ORDER))
                u_chbuffer(.memclk_i(memclk_i),
                           .channel_run_i(running),
                           .bram_uaddr_i(this_bram_uaddr),
                           .next_bram_uaddr_o(this_next_bram_uaddr),
                           .dat_i(this_channel_data),
                           .ifclk_i( ifclk_i ),
                           .bram_regce_i(this_bram_regce),
                           .bram_casdomux_i(this_bram_casdomux),
                           .bram_casdomuxen_i(this_bram_casdomuxen),
                           .bram_en_i(this_bram_en),
                           .bram_raddr_i(this_bram_raddr),
                           .dat_o(this_bram_dat_o),
                           .bram_upd_dat_i( (i==0) ? fw_dat_i : 8'h00),
                           .bram_upd_wr_i( (i==0) ? {2'b00, fw_wr_i} : 3'b000 ),
                           .bram_upd_casdimux_i( {3{1'b0}} ),
                           .cascade_in_i( cas_dinb[i] ),
                           .cascade_out_o(cas_doutb[i] ));
        end
    endgenerate        

    // flag the readout to begin
    wire readout_begin;
    // OK, here's our event header.
    // the stupidity of this cannot be overstated
    wire [31:0] header_data;
    wire header_data_valid;
    wire header_data_read;
    event_hdr_fifo u_hdr_fifo(.wr_clk(memclk_i),
                              .rd_clk(ifclk_i),
                              .rst( memclk_rst_i ),
                              .din( { event_no_i , 1'b0, trig_time_i } ),
                              .wr_en(trig_valid_i),
                              .full(),
                              .dout( header_data ),
                              .valid( header_data_valid ),
                              .rd_en( header_data_read ));
    localparam EVBITS = 3;
    localparam [EVBITS-1:0] EVIDLE = 0;
    localparam [EVBITS-1:0] HEADER_0 = 1;
    localparam [EVBITS-1:0] HEADER_1 = 2;
    localparam [EVBITS-1:0] HEADER_2 = 3;
    localparam [EVBITS-1:0] HEADER_3 = 4;
    localparam [EVBITS-1:0] DATA = 5;
    localparam [EVBITS-1:0] LAST = 6;
    reg [EVBITS-1:0] evstate = {EVBITS{1'b0}};
    reg [7:0] output_data = {8{1'b0}};
    reg       output_tlast = 0;
    reg       output_tvalid = 0;
    
    // overall sequence
    // note that we grab data on !phase, not on phase
    // and we transition on phase
    // also note that data_start_delayed is *8 CLOCKS* before
    // data becomes valid
    // clk  phase   evstate     last_data   output_data data_start_delayed  tlast
    // 0    0       EVIDLE      X           X           0                   X
    // 1    1       EVIDLE      X           X           1                   X
    // 2    0       HEADER_0    X           X           0                   X
    // 3    1       HEADER_0    X           header[0]   0                   X
    // 4    0       HEADER_1    X           header[0]   0                   X
    // 5    1       HEADER_1    X           header[1]   0                   X
    // 6    0       HEADER_2    X           header[1]   0                   X
    // 7    1       HEADER_2    X           header[2]   0                   X
    // 8    0       HEADER_3    X           header[2]   0                   X
    // 9    1       HEADER_3    data[0]     header[3]   0                   X
    // 10   0       DATA        data[0]     header[3]   0                   X
    // 11   1       DATA        data[1]     data[0]     0                   1
    // 12   0       LAST        data[1]     data[0]     0                   1
    // 13   1       LAST        X           data[1]     0                   X
    // 14   0       EVIDLE      X           data[1]     0                   X
    // etc.

    assign header_data_read = (state == LAST && dout_data_phase_i);
    
    // data_start_delayed needs to be synced up to the correct
    // phase, or else this will never work.
    always @(posedge ifclk_i) begin
        last_data_store <= last_data;
        // we capture on !phase, transition on phase
        if (ifclk_rst_i) evstate <= EVIDLE;
        else if (dout_data_phase_i) begin
            case (evstate)
                EVIDLE: if (data_start_delayed) evstate <= HEADER_0;
                HEADER_0: evstate <= HEADER_1;
                HEADER_1 : evstate <= HEADER_2;
                HEADER_2 : evstate <= HEADER_3;
                HEADER_3 : evstate <= DATA;
                DATA : if (data_tlast) evstate <= LAST;
                LAST : evstate <= EVIDLE;
            endcase
        end  
        // capture on !phase to present tvalid on phase      
        if (!dout_data_phase_i) begin
            if (evstate == HEADER_0) output_data <= header_data[31:24];
            else if (evstate == HEADER_1) output_data <= header_data[23:16];
            else if (evstate == HEADER_2) output_data <= header_data[15:8];
            else if (evstate == HEADER_3) output_data <= header_data[7:0];
            else output_data <= last_data_store;
        end
        
        if (!dout_data_phase_i) output_tlast <= (evstate == LAST);
        
        // tvalid goes high in !ifclk_phase_i if evstate != EVIDLE
        if (evstate != EVIDLE) output_tvalid <= !dout_data_phase_i;
        else output_tvalid <= 1'b0;
    end 
    
    assign dout_data_o = output_data;
    assign dout_data_valid_o= output_tvalid;
    assign dout_data_last_o = output_tlast;
        
endmodule
