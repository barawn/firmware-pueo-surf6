`timescale 1ns / 1ps
// The capture bit err detection 
module surf_sync_gen(

    );
endmodule
