`timescale 1ns / 1ps
`include "interfaces.vh"
// URAM-to-Event buffer.
// This interfaces with pueo_uram_v3+ only!
//
// We don't need a memclk_sync here -
// pueo_uram_v3+ syncs up the readout requests
// to a phase, so begin_i always occurs in phase 1.
// It's the critical timing element.
module uram_event_buffer #(parameter NCHAN = 8,
                           parameter NBIT_IN = 72,
                           parameter BEGIN_PHASE = 1,
                           parameter DOUT_LATENCY = 6)(
        input memclk_i,
        input ifclk_i,
        input begin_i,
        input [NBIT_IN*NCHAN-1:0] dat_i,
        input [NCHAN-1:0] dat_valid_i
    );
    
    localparam BEGIN_DELAY = 5;
    localparam [3:0] BEGIN_DELAY_VAL = (BEGIN_DELAY == 0) ? 0 : BEGIN_DELAY-1;
    wire begin_delayed;
    wire this_begin = (BEGIN_DELAY == 0) ? begin_i : begin_delayed;
    SRL16E u_begin_delay(.D(begin_i),
                         .CE(1'b1),
                         .CLK(memclk_i),
                         .A0(BEGIN_DELAY_VAL[0]),
                         .A1(BEGIN_DELAY_VAL[1]),
                         .A2(BEGIN_DELAY_VAL[2]),
                         .A3(BEGIN_DELAY_VAL[3]),
                         .Q(begin_delayed));
    
    // The details here are documented in the event buffer section
    // of the firmware documentation.
    // This is trickier than it first seems.
    
    // Nominally we start off by cascading the entire thing:
    // 24 total block RAMs (8 ch x 3 per channel).
    // Writing occurs at memclk speed (500 MHz), reading at ifclk speed (125 MHz)
    // So writing needs to be easy.
    
    // We write 3 addresses (24 samples) per 4 clock cycles.
    // We will ALWAYS get begin_i in phase 1.
    // Let's just consider channel 0 for the moment.
    // Suppose we register begin_i: this will then go high in phase 2.
    // We then use this signal to reset the address generation, so it's reset in phase 3.
    // The timing of a 4-address increment will always be
    // 5/6/5 6/5/6
    // This pattern is generated by the uram_event_timer.
    wire [NCHAN-1:0] channel_run;    
    // We generate a global next upper address which gets captured by ch0 and
    // forwarded.
    wire [7:0] next_bram_uaddr[NCHAN-1:0];
    // the top 3 bits are the buffer. They're Gray encoded so they can
    // hop across domains. Thankfully a 3-bit Gray counter fits in logic.

    // This is the *in progress* buffer pointer.
    // This gets incremented when the first channel finishes.
    reg [2:0] write_buffer = {3{1'b0}};
    // This is the *completed* buffer pointer. This gets incremented
    // when the last channel finishes.
    reg [2:0] complete_buffer_pointer = {3{1'b0}};
    // The reason we have 2 buffer pointers is because our control logic
    // is pipelined. We could probably just start reading out early,
    // but I'd rather be safe than sorry.
    
    // This is the upper address pointer.
    // We only pass the top 5 bits to the individual channels.
    reg [4:0] write_addr = {5{1'b0}};    
    reg [1:0] glob_memclk_phase = {2{1'b0}};
    localparam [1:0] GLOB_MEMCLK_PHASE_RESET_VAL = 3;
    wire glob_start;
    reg running = 0;
    wire increment_uaddr;
    uram_event_timer u_timer(.memclk_i(memclk_i),
                             .memclk_phase_i(!glob_memclk_phase[0]),
                             .running_i(running),
                             .start_o(glob_start),
                             .capture_o(increment_uaddr));
    always @(posedge memclk_i) begin
        if (begin_delayed) running <= 1;
        
        if (increment_uaddr) write_addr <= write_addr + 1;
        
        if (glob_start) glob_memclk_phase <= GLOB_MEMCLK_PHASE_RESET_VAL;
        else glob_memclk_phase <= glob_memclk_phase + 1;
    end                                  
    
//    assign channel_run = {NCHAN{running}};
    assign next_bram_uaddr[0] = { write_buffer, write_addr };
    generate
        genvar i;
        for (i=0;i<NCHAN;i=i+1) begin : CH
            // running delays. Looks like this should be 4*i,
            // we'll see what happens with placement and such.
            localparam RUN_DELAY = 4*i;
            // might be able to do this smarter
            if (RUN_DELAY == 0) begin : NRD
                assign channel_run[i] = running;
            end else if (RUN_DELAY < 17) begin : SRL16RD
                localparam [3:0] SRL_RUN_DLY = RUN_DELAY - 2;
                wire run_srl_delay;
                reg local_run = 0;
                SRL16E u_rundly(.D(running),
                                .CE(1'b1),
                                .CLK(memclk_i),
                                .A0(SRL_RUN_DLY[0]),
                                .A1(SRL_RUN_DLY[1]),
                                .A2(SRL_RUN_DLY[2]),
                                .A3(SRL_RUN_DLY[3]),
                                .Q(run_srl_delay));
                always @(posedge memclk_i) local_run <= run_srl_delay;
                assign channel_run[i] = local_run;                                
            end else begin : SRL32RD
                localparam [4:0] SRL_RUN_DLY = RUN_DELAY - 2;
                wire run_srl_delay;
                reg local_run = 0;
                SRLC32E u_rundly(.D(running),
                                 .CE(1'b1),
                                 .CLK(memclk_i),
                                 .A(SRL_RUN_DLY),
                                 .Q(run_srl_delay));
                always @(posedge memclk_i) local_run <= run_srl_delay;
                assign channel_run[i] = local_run;                                
            end            
            
            // this isn't *actually* synced up to memclk_sync_i:
            // it relies on the fact that channel_start is always
            // synced up because the readout sequence is.
            
            // note that our memclk phase goes 0/1/3/2 !!!
            // this is why we called it phis in the doc!
            // this is because the muxing happens A/B/B/A
            // so we can just use a single bit for that guy
            
            // reset memclk phase to this. this is actually phase 3
            localparam MEMCLK_PHASE_RESET_VAL = 0;
            // don't increment in this phase. this is actually phase 1
            localparam MEMCLK_PHASE_NO_INCREMENT = 2;
            // delay the laddr reset by this amount
            localparam LADDR_RESET_DELAY = 1;
            // select this bit from the memclk_phase to do the muxing
            localparam MEMCLK_PHASE_MUX_BIT = 1;
            // b/c of the way the muxing AND timer work,
            // we need a sequence of
            // 0 1  = 1
            // 1 0  = 2
            // 1 1  = 3
            // 0 0  = 0
            // which is just an offset count, so cool
            reg [1:0] memclk_phase = {2{1'b0}};
            reg [7:0] bram_uaddr = {8{1'b0}};
            reg [1:0] bram_laddr = {2{1'b0}};
            if (i != NCHAN-1) begin : NL
                assign next_bram_uaddr[i+1] = bram_uaddr;
            end
            wire uaddr_capture;
            wire start;
            wire reset_laddr;
            if (LADDR_RESET_DELAY == 0) begin : ND
                assign reset_laddr = start;
            end else if (LADDR_RESET_DELAY == 1) begin : RD
                reg start_rereg = 0;
                always @(posedge memclk_i) begin : DL
                    start_rereg <= start;
                end
                assign reset_laddr = start_rereg;
            end else begin : SRLD
                localparam [3:0] SRL_LADDR_DELAY_VAL = LADDR_RESET_DELAY - 1;
                SRL16E u_delay_reset(.D(start),
                                     .CE(1'b1),
                                     .CLK(memclk_i),
                                     .A0(SRL_LADDR_DELAY_VAL[0]),
                                     .A1(SRL_LADDR_DELAY_VAL[1]),
                                     .A2(SRL_LADDR_DELAY_VAL[2]),
                                     .A3(SRL_LADDR_DELAY_VAL[3]),
                                     .Q(reset_laddr));
            end
            uram_event_timer u_timer(.memclk_i(memclk_i),
                                     .memclk_phase_i(memclk_phase[0]),
                                     .running_i(channel_run[i]),
                                     .start_o(start),
                                     .capture_o(uaddr_capture));
            // ok: when start occurs that syncs us                               
            always @(posedge memclk_i) begin
                if (start) begin
                    memclk_phase <= MEMCLK_PHASE_RESET_VAL;
                end else memclk_phase <= memclk_phase + 1;
                if (reset_laddr) 
                    bram_laddr <= 2'b00;
                else if (memclk_phase != MEMCLK_PHASE_NO_INCREMENT) 
                    bram_laddr <= bram_laddr + 1;
                
                if (uaddr_capture) bram_uaddr <= next_bram_uaddr[i];                
            end                                     
        end
    endgenerate        
        
endmodule
